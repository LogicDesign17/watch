`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:10:13 06/13/2015 
// Design Name: 
// Module Name:    clock 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module clock(
    input up,
    input down,
    input left,
    input right,
    input enter,
    input esc,
    input clk,
    output [0:0] out,
    output norm,
    output [6:0] year,
    output [6:0] month,
    output [6:0] day
    );


endmodule
